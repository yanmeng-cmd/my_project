module(
    
);

endmodule